module f1_fsm(
    input   logic       clk,
    input   logic       rst,
    input   logic       en,
    input   logic       trigger,
    output  logic       cmd_seq,
    output  logic       cmd_delay,
    output  logic [7:0] data_out
);
    typedef enum  {S0, S1, S2, S3, S4, S5, S6, S7, S8} light_states;
    light_states current_state, next_state;

    always_ff @ (posedge clk)
        if (rst) current_state <= S0;
        else if (trigger & current_state==S0) current_state <= next_state;
        else if (en & current_state!=S0) current_state <= next_state;

    always_comb
        case (current_state)
            S0:     next_state = S1;
            S1:     next_state = S2;
            S2:     next_state = S3;
            S3:     next_state = S4;
            S4:     next_state = S5;
            S5:     next_state = S6;
            S6:     next_state = S7;
            S7:     next_state = S8;
            S8:     next_state = S0;
            default: next_state = S0;
        endcase

    always_comb
        case (current_state)
            S0:     data_out = 8'b0;
            S1:     data_out = 8'b1;
            S2:     data_out = 8'b11;
            S3:     data_out = 8'b111;
            S4:     data_out = 8'b1_111;
            S5:     data_out = 8'b11_111;
            S6:     data_out = 8'b111_111;
            S7:     data_out = 8'b1_111_111;
            S8:     data_out = 8'b11_111_111;
            default: data_out = 8'b0;
        endcase

    always_comb //can the syntax here be simplified? Or does this look the neatest?
        if (current_state == S8) cmd_seq = 0;
        else cmd_seq = 1;

    always_comb 
        if (current_state == S8) cmd_delay = 1;
        else cmd_delay = 0;
        
endmodule
